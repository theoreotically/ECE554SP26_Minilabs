module spart_tx(
  input clk,
  input rst,
  input enable,
  input shift_enable,
  input [7:0] txd,
  output reg tbr
);

endmodule