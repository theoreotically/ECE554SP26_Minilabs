module bus_interface(
  input        iocs,
  input        iorw,
  input        rda,
  input        tbr,
  input  [1:0] ioaddr,
  input  [7:0] rxd,
  inout  [7:0] databus,
  output [7:0] txd
);


endmodule