module spart_rx(
  input clk,
  input rst,
  input enable,
  input shift_enable,
  input [7:0] rx_bus,
  input rxd,
  output reg rda
);

endmodule