module spart_tx(
  input clk,
  input rst,
  input enable,
  input [1:0] ioaddr,
  input [7:0] txd,
  output reg tbr
);

endmodule