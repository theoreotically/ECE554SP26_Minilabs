module spart_rx(
  input clk,
  input rst,
  input enable,
  input [1:0] ioaddr,
  input rxd,
  output reg rda
);

endmodule